.SUBCKT C1206C105K1RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.239199355244637
R2 2 5 1.13999998569489
R3 1 6 1000000000
L1 1 2 3.63599983455032E-11
L2 2 3 6.90839968564561E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 7.20000028610229E-13
.param a=34 b=0.085 c=0.9
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS