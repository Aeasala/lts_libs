.SUBCKT C0805C105K3RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.0147161344527187
R2 2 5 0.509999990463257
R3 1 6 1000000000
L1 1 2 1.39999997705864E-11
L2 2 3 2.65999995641142E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 6.38000011444092E-12
.param a=15.8 b=0.23 c=0.69
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS