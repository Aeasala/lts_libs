.SUBCKT C1206C105K5RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 1.964628827571869
R2 2 5 2.54999995231628
R3 1 6 1000000000
L1 1 2 3.34999999962449E-11
L2 2 3 6.36499999928652E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 1.67999994754791E-12
.param a=22.4 b=0.16 c=0.755
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS