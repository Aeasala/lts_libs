.SUBCKT C0603C102K1RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 235.022201538086
R2 2 5 29.1999988555908
R3 1 6 99999997952
L1 1 2 1.71499994761071E-11
L2 2 3 3.25849990046034E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 2.04999995231628E-12
.param a=96 b=0.038 c=0.25
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS