.SUBCKT C0603C103K5RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.603802841318428
R2 2 5 7.18000030517578
R3 1 6 99999997952
L1 1 2 1.3500001116995E-11
L2 2 3 2.56500021222905E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 2.04999995231628E-12
.param a=50 b=0.07 c=0.239
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS