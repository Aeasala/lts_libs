.SUBCKT C1206X106K3RALTU_4x 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.912196695804596
R2 2 5 0.202500000596046
R3 1 6 25000000
L1 1 2 9.25000007145904E-12
L2 2 3 1.75750001357722E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 2.40000009536743E-12
.param a=7.6 b=0.33 c=0.92
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS