**********************************************************
*
* BC807-40
*
* Nexperia
*
* General purpose PNP transistor
* IC   = 500 mA
* VCEO = 45 V 
* hFE  = 250 - 600 @ 1V/100mA
* 
*
*
*
* Package pinning does not match Spice model pinning.
* Package: SOT 23
* 
* Package Pin 1: Base
* Package Pin 2: Emitter
* Package Pin 3: Collector
* 
*
* Extraction date (week/year): 49/2018
* Spicemodel includes temperature dependency
*
**********************************************************
*#
*
* Diode D1, Transistor Q2 and resistor RQ 
* are dedicated to improve modeling of quasi
* saturation area and reverse mode operation
* and do not reflect physical devices.
* 
.SUBCKT BC807-40 C B E
Q1 C B E Transistor 0.8544
Q2 11 B E Transistor 0.1456
RQ 11 C 19.24
*
.MODEL Transistor PNP
+ IS = 1.132E-013
+ NF = 0.9578
+ ISE = 3.045E-014
+ NE = 1.511
+ BF = 535
+ IKF = 0.2819
+ VAF = 20.46
+ NR = 0.9562
+ ISC = 3.16E-015
+ NC = 1.183
+ BR = 32
+ IKR = 0.1546
+ VAR = 12.16
+ RB = 30
+ IRB = 0.00055
+ RBM = 1.31
+ RE = 0.2017
+ RC = 0.1259
+ XTB = 1.974
+ EG = 1.11
+ XTI = 10.69
+ CJE = 4.948E-011
+ VJE = 0.6553
+ MJE = 0.3474
+ TF = 8.604E-010
+ XTF = 1.859
+ VTF = 3.813
+ ITF = 0.4203
+ PTF = 0
+ CJC = 1.786E-011
+ VJC = 0.5376
+ MJC = 0.4005
+ XCJC = 0.459
+ TR = 4.5E-008
+ CJS = 0
+ VJS = 0.75
+ MJS = 0.333
+ FC = 0.82
+ Tnom = 25
.ENDS
*