.SUBCKT C1210C106K3RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.00465048101649132
R2 2 5 0.430099993944168
R3 1 6 100000000
L1 1 2 4.49999981722016E-11
L2 2 3 8.5499996527183E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 3.25E-12
.param a=15.8 b=0.23 c=0.69
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS
