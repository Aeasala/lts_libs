.SUBCKT C0805X475K4RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 8.76356601715088
R2 2 5 1.27999997138977
R3 1 6 212800000
L1 1 2 2.33000008176276E-11
L2 2 3 4.42700015534925E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 4.03999996185303E-12
.param a=6.1 b=0.483 c=0.847
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS