.SUBCKT C1206X106K3RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.0437875837087631
R2 2 5 0.810000002384186
R3 1 6 100000000
L1 1 2 3.70000002858362E-11
L2 2 3 7.03000005430887E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 6.00000023841858E-13
.param a=7.6 b=0.33 c=0.92
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS