.SUBCKT C1206C105K3RALTU 1 6
*Temp = 25°C, Bias = 0VDC, Center Frequency = 100 Hz
*KEMET Model RLC Cerm
R1 3 4 0.260924905538559
R2 2 5 1.24000000953674
R3 1 6 1000000000
L1 1 2 3.29999999548747E-11
L2 2 3 6.26999999142619E-10
B1 4 6 I={cap*mlcc(a,b,c,abs(V(4,6)))*ddt(V(4,6))}
C2 5 6 2.04999995231628E-12
.param a=19.57 b=0.217 c=0.494
.func mlcc(a,b,c,x) {(1-(c*(0.5*(cosh(0.5*a*b)**-1)*sinh(0.5*b*x)*(cosh(0.5*b*(a-x))**-1))))}
.backanno
.end
.ENDS